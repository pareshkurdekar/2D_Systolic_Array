module corelet (clk, l0_in, l0_rd, l0_wr, reset);
  
  parameter row  = 8;
  parameter bw = 4;
  parameter col = 8; 
 
  
  input  clk;
  input [bw*col-1:0] l0_in;
  input l0_rd;
  input l0_wr;
  input reset;

  wire l0_ready;
  wire l0_full;
  reg l0_wr_q;
  wire  [row*bw-1:0] l0_out;
  
  ////////////// L0 Instance /////////////////////

    l0 #(.bw(bw)) l0_instance 
  (
        .clk(clk),
        .in(l0_in), 
        .out(l0_out), 
        .rd(l0_rd),
        .wr(l0_wr_q), 
        .o_full(l0_full), 
        .reset(reset), 
        .o_ready(l0_ready)
  );
 //////////////////////////////////////////////////////




 //////////////// IFIFO Instance ///////////////////////


 //////////////////////////////////////////////////////




 //////////////// Mac Array Instance ///////////////////


 /////////////////////////////////////////////////////



 //////////////// Ofifo Instance ///////////////////////


//////////////////////////////////////////////////////////



/////////////////////// SFP ///////////////////////////////

//////////////////////////////////////////////////////////



  always @(posedge clk)
  begin
     l0_wr_q <= l0_wr;
  end

endmodule